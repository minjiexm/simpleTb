
import uvm_pkg::*;

`include "uvm_macros.svh"
`include "apb_agent_pkg.sv"
`include "apb_test.svh"
