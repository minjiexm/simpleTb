
`include "apb_if.svh"


package apb_agent_pkg;

import uvm_pkg::*;

`include "apb_rw.svh"
`include "apb_sequences.svh"
`include "apb_driver_seq_mon.svh"
`include "apb_agent_env_config.svh"

endpackage
