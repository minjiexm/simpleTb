//
//----------------------------------------------------------------------
//   Copyright 2019 Veri5.org
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----------------------------------------------------------------------

`ifndef NETWORK_PKG_SV
`define NETWORK_PKG_SV

`include "amiq_eth_pkg.sv"

package network_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "uvme_macros.svh"
  import uvme_pkg::*;

  import amiq_eth_pkg::*;

  `include "network_macros.svh"

  `include "network_component.svh"
  `include "network_address.svh"
  `include "network_host.svh"
  `include "network_port.svh"
  `include "network_switch.svh"
  `include "network_switch_driver.svh"

endpackage : network_pkg

`endif

