//-----------------------------------------------------------------------------
//   Copyright 2019 Veri5.org
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//-----------------------------------------------------------------------------

`ifndef UVME_MACROS_SVH
`define UVME_MACROS_SVH

//
//  Include sub modules' defines
//
`include "agent/uvme_agent_defines.svh"
`include "analysis/uvme_analysis_defines.svh"
`include "args/uvme_args_defines.svh"
`include "checker/uvme_checker_defines.svh"
`include "common/uvme_common_defines.svh"
`include "event/uvme_event_pool_defines.svh"
`include "layer/uvme_layer_defines.svh"
`include "log/uvme_log_defines.svh"
`include "transaction/uvme_transaction_defines.svh"

`endif  // UVME_MACROS_SVH
